module Mux_k_to_1 
#(parameter K = 4 ,
parameter  SIZE = 16;)
(
    [SIZE - 1:0] input [0:K-1] in,
    sel,
    

);
    
endmodule