module controller(
    input clk,
    input start,
    input count_done1,
    input count_done2,
    input carry2,
    input carry3,
    input carry4,
);
    


endmodule