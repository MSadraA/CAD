module inv_mod(
    input a,
    output b
);

    assign b = (~a);

endmodule