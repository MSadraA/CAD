module controller(
    input clk,
    input start,
    input count_done1,
    input count_done2,
    
);

endmodule