module IfMapSP #(
    parameter DATA_WIDTH = 16,
    parameter SIZE = 16
) (
    input clk, 
    input rst,
    input[DATA_WIDTH - 1 : 0] din,
    input $clog2()
);
    
endmodule